ddd

dddxxxxxd
